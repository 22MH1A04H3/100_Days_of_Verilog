module name_tb;
reg [5:0]a;
wire y;
name uut(.a(a),.y(y));
initial
begin
a=6'b111111;//D
#5;
a=6'b100001;
#5;
a=6'b100001;
#5;
a=6'b011110;
#5;
a=6'b000000;
#5;
a=6'b111111;//A
#5;
a=6'b001001;
#5;

a=6'b001001;
#5;

a=6'b111111;
#5;
a=6'b000000;
#5;
a=6'b110111;//s
#5;
a=6'b100101;
#5;
a=6'b100101;
#5;
a=6'b111101;
#5;
a=6'b000000;
#5;

a=6'b111111;//u
#5;

a=6'b100000;
#5;

a=6'b100000;
#5;
a=6'b111111;
#5;
a=6'b000000;
#5;
a=6'b111111;//k
#5;
a=6'b000100;
#5;
a=6'b001010;
#5;
a=6'b110001;
#5;
a=6'b000000;
#5;
a=6'b111111;//o
#5;
a=6'b100001;
#5;
a=6'b100001;
#5;
a=6'b111111;
#5;
a=6'b000000;
#5;
a=6'b111111;//D
#5;
a=6'b100001;
#5;
a=6'b100001;
#5;
a=6'b011110;
#5;
a=6'b000000;
#5;
a=6'b111111;//A
#5;
a=6'b001001;
#5;

a=6'b001001;
#5;

a=6'b111111;
#5;
a=6'b000000;
#5;

$finish();
end
endmodule
