//verilog HDL to generate clk with 100MHZ
module clk_gen(
input clk);
endmodule
